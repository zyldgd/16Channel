/*
 * file   : LTC220X_data_sampling.v
 * author : zyl
 * date   : 2018-8-22
 * addr   : whu.edu.ionosphereLab
 */

module LTC220X_data_sampling(
input   

);

endmodule 
//end LTC220X_data_sampling